--------------------------------------------------------------------------
--
-- SysConCharRom
--
-- Character ROM for SysCon's video controller
-- (128 characters with box draw characters in < 32)
-- 
-- Copyright (C) 2019 Topten Software.  All Rights Reserved.
--
--------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;
use std.textio.all;
use ieee.std_logic_textio.all;

entity SysConCharRom is
port
(
	i_clock : in std_logic;
	i_addr : in std_logic_vector(10 downto 0);
	o_dout : out std_logic_vector(7 downto 0)
);
end SysConCharRom;

--xilt:nowarn:Signal 'ram', unconnected in block 'SysConCharRom', is tied to its initial value.
 
architecture behavior of SysConCharRom is 
	type mem_type is array(0 to 2047) of std_logic_vector(7 downto 0);
	signal ram : mem_type := (
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"ff", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"f0", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", 
x"10", x"10", x"10", x"10", x"10", x"1f", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"10", x"10", x"10", x"10", x"10", x"f0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"1f", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", 
x"10", x"10", x"10", x"10", x"10", x"ff", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"ff", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", 
x"10", x"10", x"10", x"10", x"10", x"1f", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", 
x"10", x"10", x"10", x"10", x"10", x"f0", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", 
x"10", x"10", x"10", x"10", x"10", x"ff", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", 
x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"00", x"00", x"00", 
x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"00", x"00", x"00", x"00", 
x"0f", x"0f", x"0f", x"0f", x"0f", x"0f", x"0f", x"0f", x"0f", x"0f", x"0f", x"0f", x"00", x"00", x"00", x"00", 
x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"0f", x"0f", x"0f", x"0f", x"0f", x"0f", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"0f", x"0f", x"0f", x"0f", x"0f", x"0f", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"00", x"00", x"00", x"00", 
x"00", x"00", x"3c", x"3c", x"3c", x"3c", x"3c", x"3c", x"3c", x"3c", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"10", x"10", x"38", x"38", x"7c", x"7c", x"fe", x"fe", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"fe", x"fe", x"7c", x"7c", x"38", x"38", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"80", x"c0", x"e0", x"f8", x"fe", x"f8", x"e0", x"c0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"02", x"06", x"0e", x"3e", x"fe", x"3e", x"0e", x"06", x"02", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"08", x"1c", x"2a", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"08", x"08", x"2a", x"1c", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"10", x"08", x"7c", x"08", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"08", x"10", x"3e", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"55", x"aa", x"55", x"aa", x"55", x"aa", x"55", x"aa", x"55", x"aa", x"55", x"aa", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"10", x"10", x"10", x"10", x"10", x"00", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"28", x"28", x"28", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"28", x"28", x"7c", x"28", x"7c", x"28", x"28", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"10", x"3c", x"50", x"38", x"14", x"78", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"60", x"64", x"08", x"10", x"20", x"4c", x"0c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"20", x"50", x"50", x"20", x"54", x"48", x"34", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"30", x"30", x"20", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"08", x"10", x"20", x"20", x"20", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"20", x"10", x"08", x"08", x"08", x"10", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"10", x"54", x"38", x"7c", x"38", x"54", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"10", x"10", x"7c", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"20", x"40", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"7c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"04", x"08", x"10", x"20", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"44", x"4c", x"54", x"64", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"10", x"30", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"44", x"04", x"38", x"40", x"40", x"7c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"44", x"04", x"18", x"04", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"08", x"18", x"28", x"48", x"7c", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"7c", x"40", x"38", x"04", x"04", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"18", x"20", x"40", x"78", x"44", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"7c", x"04", x"08", x"10", x"20", x"40", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"44", x"44", x"38", x"44", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"44", x"44", x"3c", x"04", x"08", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"30", x"30", x"00", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"30", x"30", x"00", x"30", x"30", x"20", x"40", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"08", x"10", x"20", x"40", x"20", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"7c", x"00", x"7c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"20", x"10", x"08", x"04", x"08", x"10", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"44", x"04", x"08", x"10", x"00", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"44", x"04", x"34", x"54", x"54", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"10", x"28", x"44", x"44", x"7c", x"44", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"78", x"24", x"24", x"38", x"24", x"24", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"44", x"40", x"40", x"40", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"78", x"24", x"24", x"24", x"24", x"24", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"7c", x"40", x"40", x"70", x"40", x"40", x"7c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"7c", x"40", x"40", x"70", x"40", x"40", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"3c", x"40", x"40", x"4c", x"44", x"44", x"3c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"44", x"44", x"44", x"7c", x"44", x"44", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"10", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"04", x"04", x"04", x"04", x"04", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"44", x"48", x"50", x"60", x"50", x"48", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"40", x"40", x"40", x"40", x"40", x"40", x"7c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"44", x"6c", x"54", x"54", x"44", x"44", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"44", x"64", x"54", x"4c", x"44", x"44", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"44", x"44", x"44", x"44", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"78", x"44", x"44", x"78", x"40", x"40", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"44", x"44", x"44", x"54", x"48", x"34", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"78", x"44", x"44", x"78", x"50", x"48", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"44", x"40", x"38", x"04", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"7c", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"44", x"44", x"44", x"44", x"44", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"44", x"44", x"44", x"28", x"28", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"44", x"44", x"44", x"44", x"54", x"6c", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"44", x"44", x"28", x"10", x"28", x"44", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"44", x"44", x"28", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"7c", x"04", x"08", x"10", x"20", x"40", x"7c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"20", x"20", x"20", x"20", x"20", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"40", x"20", x"10", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"38", x"08", x"08", x"08", x"08", x"08", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"10", x"28", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"18", x"18", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"38", x"04", x"3c", x"44", x"3c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"40", x"40", x"58", x"64", x"44", x"64", x"58", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"38", x"44", x"40", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"04", x"04", x"34", x"4c", x"44", x"4c", x"34", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"38", x"44", x"7c", x"40", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"08", x"14", x"10", x"38", x"10", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"34", x"4c", x"4c", x"34", x"04", x"44", x"38", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"40", x"40", x"58", x"64", x"44", x"44", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"10", x"00", x"30", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"04", x"00", x"04", x"04", x"04", x"04", x"44", x"38", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"40", x"40", x"48", x"50", x"60", x"50", x"48", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"30", x"10", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"68", x"54", x"54", x"54", x"54", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"58", x"64", x"44", x"44", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"38", x"44", x"44", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"58", x"64", x"44", x"64", x"58", x"40", x"40", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"34", x"4c", x"44", x"4c", x"34", x"04", x"04", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"58", x"64", x"40", x"40", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"3c", x"40", x"38", x"04", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"10", x"10", x"7c", x"10", x"10", x"14", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"44", x"44", x"44", x"4c", x"34", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"44", x"44", x"44", x"28", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"44", x"44", x"54", x"54", x"28", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"44", x"28", x"10", x"28", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"44", x"44", x"44", x"3c", x"04", x"44", x"38", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"7c", x"08", x"10", x"20", x"7c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"08", x"10", x"10", x"20", x"10", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"10", x"10", x"10", x"00", x"10", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"20", x"10", x"10", x"08", x"10", x"10", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"20", x"54", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"28", x"54", x"28", x"54", x"28", x"54", x"28", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
);
begin

	process (i_clock)
	begin
		if rising_edge(i_clock) then

			o_dout <= ram(to_integer(unsigned(i_addr)));

		end if;
	end process;
end;
